//Control store controls all signals

module LC3_controlstore(
    //This module stores the microinstrustions
    input clk,
    
);
endmodule